-- --------------------------------------------------------------------
--
-- Future copywrite / licensing information?
--
-- ...
--
-- ...
--
--   Title     :  Package(s) Names
--             :  (PACKAGE_NAME package declaration)
--             :
--   Library   :  library info
--             :
--   Developers:  Davis Rash
--             :
--   Purpose   :  purpose!
--             :
--   Limitation:  very limited!
--             :
--   Note      : more notes
--             :
-- --------------------------------------------------------------------
-- $Revision: 0 $
-- $Date: YYYY-MM-DD HH:MM:SS +XXXX (DOW, DD Mon YYYY) $
-- --------------------------------------------------------------------

-- use STD.TEXTIO.all;
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package body vectors is

end package body vectors;
